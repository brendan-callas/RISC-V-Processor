import rv32i_types::*;

module datapath
(

);



endmodule : datapath